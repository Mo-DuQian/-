`include "lib/defines.vh"
module EX(
    input wire clk,
    input wire rst,
    // input wire flush,
    input wire [`StallBus-1:0] stall,

    input wire [`ID_TO_EX_WD-1:0] id_to_ex_bus,

    output wire [`EX_TO_MEM_WD-1:0] ex_to_mem_bus,

    output wire data_sram_en,
    output wire [3:0] data_sram_wen,
    output wire [31:0] data_sram_addr,
    output wire [31:0] data_sram_wdata,
    
    //���ex�������
    output wire [4:0] cf_ex_addr,
    output wire [31:0] cf_ex_data,
    output wire cf_ex_we,
    
    output wire [5:0] ex_opcode,
    
    output wire cf_ex_we_hi,
    output wire cf_ex_we_lo,
    output wire [31:0] cf_ex_hi,
    output wire [31:0] cf_ex_lo,
    
    output wire stallreq_for_ex
);

    reg [`ID_TO_EX_WD-1:0] id_to_ex_bus_r;

    always @ (posedge clk) begin
        if (rst) begin
            id_to_ex_bus_r <= `ID_TO_EX_WD'b0;
        end
        // else if (flush) begin
        //     id_to_ex_bus_r <= `ID_TO_EX_WD'b0;
        // end
        else if (stall[2]==`Stop && stall[3]==`NoStop) begin
            id_to_ex_bus_r <= `ID_TO_EX_WD'b0;
        end
        else if (stall[2]==`NoStop) begin
            id_to_ex_bus_r <= id_to_ex_bus;
        end
    end

    wire [31:0] ex_pc, inst;
    wire [11:0] alu_op;
    wire [2:0] sel_alu_src1;
    wire [6:0] sel_alu_src2;
    wire data_ram_en;
    wire [3:0] data_ram_wen;
    wire rf_we;
    wire [4:0] rf_waddr;
    wire sel_rf_res;
    wire [31:0] rf_rdata1, rf_rdata2;
    reg is_in_delayslot; //�����ô����
    
    wire ex_we_hi;
    wire ex_we_lo;
    wire [31:0] ex_hi_i,ex_hi;
    wire [31:0] ex_lo_i,ex_lo;
    
    wire inst_div, inst_divu;
    wire inst_mult,inst_multu;
    wire inst_lb,inst_lbu,inst_lh,inst_lhu,inst_sb,inst_sh;

    assign {
        inst_lb,
        inst_lbu,
        inst_lh,
        inst_lhu,
        inst_sb,
        inst_sh,
        inst_mult,
        inst_multu,
        inst_div,
        inst_divu,
        ex_we_hi,
        ex_we_lo,
        ex_hi_i,
        ex_lo_i,
        ex_pc,          // 148:117
        inst,           // 116:85
        alu_op,         // 84:83
        sel_alu_src1,   // 82:80 //��չ�˼�λ
        sel_alu_src2,   // 79:76
        data_ram_en,    // 75
        data_ram_wen,   // 74:71
        rf_we,          // 70
        rf_waddr,       // 69:65
        sel_rf_res,     // 64
        rf_rdata1,         // 63:32
        rf_rdata2          // 31:0
    } = id_to_ex_bus_r;
    
    assign ex_opcode = inst[31:26];
    wire [31:0] imm_sign_extend, imm_zero_extend, sa_zero_extend;
    assign imm_sign_extend = {{16{inst[15]}},inst[15:0]};
    assign imm_zero_extend = {16'b0, inst[15:0]};
    assign sa_zero_extend = {27'b0,inst[10:6]};

    wire [31:0] alu_src1, alu_src2;
    wire [31:0] alu_result, ex_result;
    //assign data_sram_en = data_ram_en;
    //assign data_sram_wen = data_ram_wen;
    //assign data_sram_addr = ex_result;
    //assign data_sram_wdata = rf_rdata2;

    assign alu_src1 = sel_alu_src1[1] ? ex_pc :
                      sel_alu_src1[2] ? sa_zero_extend : 
                      rf_rdata1;

    assign alu_src2 = sel_alu_src2[1] ? imm_sign_extend :
                      sel_alu_src2[2] ? 32'd8 :
                      sel_alu_src2[3] ? imm_zero_extend : 
                      sel_alu_src2[4] ? ex_lo_i :
                      sel_alu_src2[5] ? ex_hi_i:
                      sel_alu_src2[6] ? 32'b0:
                      rf_rdata2;
    
    alu u_alu(
    	.alu_control (alu_op ),
        .alu_src1    (alu_src1    ),
        .alu_src2    (alu_src2    ),
        .alu_result  (alu_result  )
    );
    
    
    assign data_sram_en = data_ram_en;
    
    
    assign data_sram_wen =  inst_sb & alu_result[1:0] == 2'b00 ? 4'b0001:
                            inst_sb & alu_result[1:0] == 2'b01 ? 4'b0010:
                            inst_sb & alu_result[1:0] == 2'b10 ? 4'b0100:
                            inst_sb & alu_result[1:0] == 2'b11 ? 4'b1000:
                            inst_sh & alu_result[1:0] == 2'b00 ? 4'b0011:
                            inst_sh & alu_result[1:0] == 2'b10 ? 4'b1100:
                            data_ram_wen;
    assign data_sram_addr = ex_result; //������alu_result
    //assign data_sram_wdata = rf_rdata2;
//    assign data_sram_wdata = data_sram_wen==4'b0001 ? {24'b0,rf_rdata2[7:0]}:
//                             data_sram_wen==4'b0010 ? {24'b0,rf_rdata2[15:8]}:
//                             data_sram_wen==4'b0100 ? {24'b0,rf_rdata2[23:16]}:
//                             data_sram_wen==4'b1000 ? {24'b0,rf_rdata2[31:24]}:
//                             data_sram_wen==4'b0011 ? {16'b0,rf_rdata2[15:0]}:
//                             data_sram_wen==4'b1100 ? {16'b0,rf_rdata2[31:16]}:
//                             rf_rdata2;

    assign data_sram_wdata = data_sram_wen==4'b0001 ? {rf_rdata2[7:0],rf_rdata2[7:0],rf_rdata2[7:0],rf_rdata2[7:0]}:
                             data_sram_wen==4'b0010 ? {rf_rdata2[7:0],rf_rdata2[7:0],rf_rdata2[7:0],rf_rdata2[7:0]}:
                             data_sram_wen==4'b0100 ? {rf_rdata2[7:0],rf_rdata2[7:0],rf_rdata2[7:0],rf_rdata2[7:0]}:
                             data_sram_wen==4'b1000 ? {rf_rdata2[7:0],rf_rdata2[7:0],rf_rdata2[7:0],rf_rdata2[7:0]}:
                             data_sram_wen==4'b0011 ? {rf_rdata2[15:0],rf_rdata2[15:0]}:
                             data_sram_wen==4'b1100 ? {rf_rdata2[15:0],rf_rdata2[15:0]}:
                             rf_rdata2;
    
    
    // MUL part
    wire [63:0] mul_result;
    wire mul_signed; // �з��ų˷����
    assign mul_signed = inst_mult;
    

    mul u_mul(
    	.clk        (clk            ),
        .resetn     (~rst           ),
        .mul_signed (mul_signed     ),
        .ina        ( alu_src1     ), // �˷�Դ������1
        .inb        ( alu_src2     ), // �˷�Դ������2  
        .result     (mul_result     ) // �˷���� 64bit
    );

    // DIV part
    wire [63:0] div_result;
    //wire inst_div, inst_divu;
    wire div_ready_i;
    reg stallreq_for_div;
    assign stallreq_for_ex = stallreq_for_div;
    
    

    reg [31:0] div_opdata1_o;
    reg [31:0] div_opdata2_o;
    reg div_start_o;
    reg signed_div_o;

    div u_div(
    	.rst          (rst          ),
        .clk          (clk          ),
        .signed_div_i (signed_div_o ),
        .opdata1_i    (div_opdata1_o    ),
        .opdata2_i    (div_opdata2_o    ),
        .start_i      (div_start_o      ),
        .annul_i      (1'b0      ),
        .result_o     (div_result     ), // ������� 64bit
        .ready_o      (div_ready_i      )
    );

    always @ (*) begin
        if (rst) begin
            stallreq_for_div = `NoStop;
            div_opdata1_o = `ZeroWord;
            div_opdata2_o = `ZeroWord;
            div_start_o = `DivStop;
            signed_div_o = 1'b0;
        end
        else begin
            stallreq_for_div = `NoStop;
            div_opdata1_o = `ZeroWord;
            div_opdata2_o = `ZeroWord;
            div_start_o = `DivStop;
            signed_div_o = 1'b0;
            case ({inst_div,inst_divu})
                2'b10:begin
                    if (div_ready_i == `DivResultNotReady) begin
                        div_opdata1_o = rf_rdata1;
                        div_opdata2_o = rf_rdata2;
                        div_start_o = `DivStart;
                        signed_div_o = 1'b1;
                        stallreq_for_div = `Stop;
                        
                    end
                    else if (div_ready_i == `DivResultReady) begin
                        div_opdata1_o = rf_rdata1;
                        div_opdata2_o = rf_rdata2;
                        div_start_o = `DivStop;
                        signed_div_o = 1'b1;
                        stallreq_for_div = `NoStop;
                    end
                    else begin
                        div_opdata1_o = `ZeroWord;
                        div_opdata2_o = `ZeroWord;
                        div_start_o = `DivStop;
                        signed_div_o = 1'b0;
                        stallreq_for_div = `NoStop;
                    end
                end
                2'b01:begin
                    if (div_ready_i == `DivResultNotReady) begin
                        div_opdata1_o = rf_rdata1;
                        div_opdata2_o = rf_rdata2;
                        div_start_o = `DivStart;
                        signed_div_o = 1'b0;
                        stallreq_for_div = `Stop;
                    end
                    else if (div_ready_i == `DivResultReady) begin
                        div_opdata1_o = rf_rdata1;
                        div_opdata2_o = rf_rdata2;
                        div_start_o = `DivStop;
                        signed_div_o = 1'b0;
                        stallreq_for_div = `NoStop;
                    end
                    else begin
                        div_opdata1_o = `ZeroWord;
                        div_opdata2_o = `ZeroWord;
                        div_start_o = `DivStop;
                        signed_div_o = 1'b0;
                        stallreq_for_div = `NoStop;
                    end
                end
                default:begin
                end
            endcase
        end
    end

    // mul_result �� div_result ����ֱ��ʹ��
    
    //assign stallreq_for_ex = stallreq_for_div;
    
    assign ex_result = alu_result;  
    
    assign ex_hi=ex_we_hi & (inst_div| inst_divu)? div_result[63:32] :
                 ex_we_hi & (inst_mult| inst_multu)? mul_result[63:32] :
                 ex_we_hi ? alu_result :   
                 ex_hi_i; 
    assign ex_lo=ex_we_lo & (inst_div | inst_divu) ? div_result[31:0] :
                 ex_we_lo & (inst_mult | inst_multu) ? mul_result[31:0] :
                 ex_we_lo ? alu_result :
                 ex_lo_i;
    
    assign cf_ex_we = rf_we;
    assign cf_ex_addr = rf_waddr;
    assign cf_ex_data = ex_result;
    
    assign cf_ex_we_hi=ex_we_hi;//��������Ҫ���ж�
    assign cf_ex_we_lo=ex_we_lo;
    assign cf_ex_hi = ex_hi;
    assign cf_ex_lo = ex_lo;
    
    
                    
     

    assign ex_to_mem_bus = {
        inst_lb,
        inst_lbu,
        inst_lh,
        inst_lhu,
        ex_we_hi,
        ex_we_lo,
        ex_hi,
        ex_lo,
        ex_pc,          // 75:44
        data_ram_en,    // 43
        data_ram_wen,   // 42:39
        sel_rf_res,     // 38
        rf_we,          // 37
        rf_waddr,       // 36:32
        ex_result       // 31:0
    };
    
    
    
endmodule